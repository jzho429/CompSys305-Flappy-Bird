-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.0 Build 156 04/24/2013 SJ Full Version
-- Created on Tue May 25 16:49:14 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY flappyBirdState IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        dead : IN STD_LOGIC := '0';
        mouseLeft : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        mouseRight : IN STD_LOGIC := '0';
        mouseRow : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
        mouseCol : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
        stateOut : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
    );
END flappyBirdState;

ARCHITECTURE BEHAVIOR OF flappyBirdState IS
    TYPE type_fstate IS (menu,idleT,idle1,idle2,idle3,lvlT,lvl1,lvl2,lvl3,death);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,dead,mouseLeft,mouseRight,mouseRow,mouseCol)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= menu;
            stateOut <= "000";
        ELSE
            stateOut <= "000";
            CASE fstate IS
                WHEN menu =>
                    IF ((((mouseLeft(1 DOWNTO 0) = "01") AND ((mouseRow(9 DOWNTO 0) >= "0011110000") AND (mouseRow(9 DOWNTO 0) < "0100001100"))) AND ((mouseCol(9 DOWNTO 0) >= "0100011000") AND (mouseCol(9 DOWNTO 0) < "0101101000")))) THEN
                        reg_fstate <= idleT;
                    ELSIF ((((mouseLeft(1 DOWNTO 0) = "01") AND ((mouseRow(9 DOWNTO 0) >= "0100011100") AND (mouseRow(9 DOWNTO 0) < "0100110110"))) AND ((mouseCol(9 DOWNTO 0) >= "0100011000") AND (mouseCol(9 DOWNTO 0) < "0101101000")))) THEN
                        reg_fstate <= idle1;
                    ELSIF ((((mouseLeft(1 DOWNTO 0) = "01") AND ((mouseRow(9 DOWNTO 0) >= "0101000100") AND (mouseRow(9 DOWNTO 0) < "0101100000"))) AND ((mouseCol(9 DOWNTO 0) >= "0100011000") AND (mouseCol(9 DOWNTO 0) < "0101101000")))) THEN
                        reg_fstate <= idle2;
                    ELSIF ((((mouseLeft(1 DOWNTO 0) = "01") AND ((mouseRow(9 DOWNTO 0) >= "0101101110") AND (mouseRow(9 DOWNTO 0) < "0110001010"))) AND ((mouseCol(9 DOWNTO 0) >= "0100011000") AND (mouseCol(9 DOWNTO 0) < "0101101000")))) THEN
                        reg_fstate <= idle3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= menu;
                    END IF;

                    stateOut <= "000";
                WHEN idleT =>
                    IF ((mouseLeft(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= lvlT;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= idleT;
                    END IF;

                    stateOut <= "001";
                WHEN idle1 =>
                    IF ((mouseLeft(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= lvl1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= idle1;
                    END IF;

                    stateOut <= "001";
                WHEN idle2 =>
                    IF ((mouseLeft(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= lvl2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= idle2;
                    END IF;

                    stateOut <= "001";
                WHEN idle3 =>
                    IF ((mouseLeft(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= lvl3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= idle3;
                    END IF;

                    stateOut <= "001";
                WHEN lvlT =>
                    IF ((mouseRight = '1')) THEN
                        reg_fstate <= menu;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= lvlT;
                    END IF;

                    stateOut <= "010";
                WHEN lvl1 =>
                    IF ((dead = '1')) THEN
                        reg_fstate <= death;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= lvl1;
                    END IF;

                    stateOut <= "011";
                WHEN lvl2 =>
                    IF ((dead = '1')) THEN
                        reg_fstate <= death;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= lvl2;
                    END IF;

                    stateOut <= "100";
                WHEN lvl3 =>
                    IF ((dead = '1')) THEN
                        reg_fstate <= death;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= lvl3;
                    END IF;

                    stateOut <= "101";
                WHEN death =>
                    IF ((((mouseLeft(1 DOWNTO 0) = "01") AND ((mouseRow(9 DOWNTO 0) >= "0011110000") AND (mouseRow(9 DOWNTO 0) < "0100001100"))) AND ((mouseCol(9 DOWNTO 0) >= "0100011000") AND (mouseCol(9 DOWNTO 0) < "0101101000")))) THEN
                        reg_fstate <= menu;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= death;
                    END IF;

                    stateOut <= "110";
                WHEN OTHERS => 
                    stateOut <= "XXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
